

module delay_line (input clk, input rst_n
    ,input din, output dout
    ,input [11:0] delay
);



endmodule


