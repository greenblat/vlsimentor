
module pld30 (

// programming interface, shift register style
     input prog_clk
    ,input prog_data

// functional  interface
    ,input [29:0] din
    ,output [29:0] dout
);


// put Your imagination here
// DONT SHARE YOUR DESIGN with me. I am working on it too!!!!

endmodule


