module rnd (input [7:0] sel, output reg [7:0] rndout);

always @* begin
    case (sel)
        0 : rndout = 19;
        1 : rndout = 213;
        2 : rndout = 208;
        3 : rndout = 31;
        4 : rndout = 161;
        5 : rndout = 104;
        6 : rndout = 201;
        7 : rndout = 153;
        8 : rndout = 77;
        9 : rndout = 182;
        10 : rndout = 192;
        11 : rndout = 20;
        12 : rndout = 216;
        13 : rndout = 121;
        14 : rndout = 44;
        15 : rndout = 225;
        16 : rndout = 94;
        17 : rndout = 203;
        18 : rndout = 211;
        19 : rndout = 36;
        20 : rndout = 23;
        21 : rndout = 24;
        22 : rndout = 165;
        23 : rndout = 216;
        24 : rndout = 54;
        25 : rndout = 113;
        26 : rndout = 133;
        27 : rndout = 25;
        28 : rndout = 247;
        29 : rndout = 175;
        30 : rndout = 200;
        31 : rndout = 214;
        32 : rndout = 230;
        33 : rndout = 194;
        34 : rndout = 31;
        35 : rndout = 174;
        36 : rndout = 81;
        37 : rndout = 148;
        38 : rndout = 176;
        39 : rndout = 237;
        40 : rndout = 102;
        41 : rndout = 221;
        42 : rndout = 103;
        43 : rndout = 246;
        44 : rndout = 130;
        45 : rndout = 252;
        46 : rndout = 68;
        47 : rndout = 157;
        48 : rndout = 197;
        49 : rndout = 116;
        50 : rndout = 49;
        51 : rndout = 167;
        52 : rndout = 75;
        53 : rndout = 112;
        54 : rndout = 180;
        55 : rndout = 193;
        56 : rndout = 126;
        57 : rndout = 91;
        58 : rndout = 221;
        59 : rndout = 217;
        60 : rndout = 255;
        61 : rndout = 193;
        62 : rndout = 218;
        63 : rndout = 144;
        64 : rndout = 152;
        65 : rndout = 193;
        66 : rndout = 167;
        67 : rndout = 214;
        68 : rndout = 122;
        69 : rndout = 0;
        70 : rndout = 80;
        71 : rndout = 30;
        72 : rndout = 195;
        73 : rndout = 10;
        74 : rndout = 78;
        75 : rndout = 98;
        76 : rndout = 25;
        77 : rndout = 107;
        78 : rndout = 83;
        79 : rndout = 91;
        80 : rndout = 210;
        81 : rndout = 222;
        82 : rndout = 6;
        83 : rndout = 178;
        84 : rndout = 69;
        85 : rndout = 195;
        86 : rndout = 134;
        87 : rndout = 85;
        88 : rndout = 211;
        89 : rndout = 77;
        90 : rndout = 49;
        91 : rndout = 248;
        92 : rndout = 68;
        93 : rndout = 105;
        94 : rndout = 123;
        95 : rndout = 21;
        96 : rndout = 173;
        97 : rndout = 10;
        98 : rndout = 205;
        99 : rndout = 116;
        100 : rndout = 61;
        101 : rndout = 216;
        102 : rndout = 165;
        103 : rndout = 112;
        104 : rndout = 38;
        105 : rndout = 161;
        106 : rndout = 235;
        107 : rndout = 238;
        108 : rndout = 148;
        109 : rndout = 96;
        110 : rndout = 213;
        111 : rndout = 149;
        112 : rndout = 189;
        113 : rndout = 144;
        114 : rndout = 47;
        115 : rndout = 191;
        116 : rndout = 197;
        117 : rndout = 166;
        118 : rndout = 56;
        119 : rndout = 177;
        120 : rndout = 156;
        121 : rndout = 49;
        122 : rndout = 174;
        123 : rndout = 240;
        124 : rndout = 51;
        125 : rndout = 174;
        126 : rndout = 247;
        127 : rndout = 176;
        128 : rndout = 143;
        129 : rndout = 152;
        130 : rndout = 224;
        131 : rndout = 66;
        132 : rndout = 108;
        133 : rndout = 86;
        134 : rndout = 167;
        135 : rndout = 130;
        136 : rndout = 17;
        137 : rndout = 169;
        138 : rndout = 59;
        139 : rndout = 65;
        140 : rndout = 133;
        141 : rndout = 135;
        142 : rndout = 233;
        143 : rndout = 77;
        144 : rndout = 205;
        145 : rndout = 129;
        146 : rndout = 36;
        147 : rndout = 71;
        148 : rndout = 223;
        149 : rndout = 209;
        150 : rndout = 39;
        151 : rndout = 109;
        152 : rndout = 11;
        153 : rndout = 65;
        154 : rndout = 12;
        155 : rndout = 188;
        156 : rndout = 67;
        157 : rndout = 139;
        158 : rndout = 153;
        159 : rndout = 46;
        160 : rndout = 30;
        161 : rndout = 49;
        162 : rndout = 5;
        163 : rndout = 179;
        164 : rndout = 240;
        165 : rndout = 170;
        166 : rndout = 17;
        167 : rndout = 123;
        168 : rndout = 57;
        169 : rndout = 82;
        170 : rndout = 153;
        171 : rndout = 95;
        172 : rndout = 223;
        173 : rndout = 150;
        174 : rndout = 156;
        175 : rndout = 205;
        176 : rndout = 148;
        177 : rndout = 98;
        178 : rndout = 87;
        179 : rndout = 3;
        180 : rndout = 40;
        181 : rndout = 18;
        182 : rndout = 224;
        183 : rndout = 194;
        184 : rndout = 144;
        185 : rndout = 86;
        186 : rndout = 5;
        187 : rndout = 5;
        188 : rndout = 138;
        189 : rndout = 94;
        190 : rndout = 87;
        191 : rndout = 245;
        192 : rndout = 22;
        193 : rndout = 39;
        194 : rndout = 102;
        195 : rndout = 166;
        196 : rndout = 199;
        197 : rndout = 40;
        198 : rndout = 39;
        199 : rndout = 215;
        200 : rndout = 106;
        201 : rndout = 11;
        202 : rndout = 204;
        203 : rndout = 223;
        204 : rndout = 185;
        205 : rndout = 9;
        206 : rndout = 240;
        207 : rndout = 167;
        208 : rndout = 16;
        209 : rndout = 51;
        210 : rndout = 164;
        211 : rndout = 242;
        212 : rndout = 142;
        213 : rndout = 255;
        214 : rndout = 26;
        215 : rndout = 122;
        216 : rndout = 239;
        217 : rndout = 53;
        218 : rndout = 41;
        219 : rndout = 199;
        220 : rndout = 75;
        221 : rndout = 85;
        222 : rndout = 132;
        223 : rndout = 53;
        224 : rndout = 216;
        225 : rndout = 32;
        226 : rndout = 126;
        227 : rndout = 108;
        228 : rndout = 125;
        229 : rndout = 186;
        230 : rndout = 169;
        231 : rndout = 18;
        232 : rndout = 153;
        233 : rndout = 203;
        234 : rndout = 237;
        235 : rndout = 76;
        236 : rndout = 46;
        237 : rndout = 77;
        238 : rndout = 150;
        239 : rndout = 34;
        240 : rndout = 52;
        241 : rndout = 124;
        242 : rndout = 215;
        243 : rndout = 136;
        244 : rndout = 125;
        245 : rndout = 150;
        246 : rndout = 180;
        247 : rndout = 30;
        248 : rndout = 26;
        249 : rndout = 215;
        250 : rndout = 40;
        251 : rndout = 64;
        252 : rndout = 4;
        253 : rndout = 120;
        254 : rndout = 13;
        255 : rndout = 46;
        default: rndout = 0;
    endcase
end
endmodule


