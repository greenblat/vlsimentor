`define PLUG_RGF_BASEADDR    'h0
`define ADDR_CONTROL                                             'h0
`define ADDR_STATUS                                              'hc
`define ADDR_CONTROL2                                            'h10
