
module pld30 (
     input prog_clk
    ,input prog_data
    ,input [29:0] din
    ,output [29:0] dout
);


// put Your imagination here

endmodule


